library ieee;
use i